`define DRAM_CYCLE    30.4
`define ROM_CYCLE     50.2
`define SRAM_CYCLE    11.0
`define CPU_CYCLE     12.5
`define AXI_CYCLE     25.0 // 40Mhz
